/*
 ------------------------------------------------------------------------------
 -
 - FILE        : bench.v 
 - Design      : FIX Engine
 - Description : Automated testbench for design
 - Author      : Adil Sadik <sadik.adil@gmail.com, ams2378@columbia.edu> 
 -
 -----------------------------------------------------------------------------
 -
 - Created     : 03/26/2013
 - Revision    : 03/30/2013 
 -		 Included Verilog-event feature for better control 
 -		 over execution flow   
 -
 -		
 -
 -----------------------------------------------------------------------------
 -
 -  Dependency  : dut.v, init_in.txt, init_out.txt
 -  Output Log  : monitor.txt
 -   
 -  Status	: Only deals with Initiator side. 
 -		  Good (compiling and dumping waveforms in desired format)
 -  TODO	: Need to add acceptor side (should be very trivial)	  
 -   		  Need real DUT for verification (in progress)
 -   
 -  Instruction : For simulation, run "sh runsim.sh" from command line
 -		  Sim log saved in "transcript"		
 -		  Run "nuke.sh" to clean the dir
 -		  
 - needtodefine: file: logon, heartbeat
 -	  	 states: connected, logonsent, waiting_for_connection, heartbeatsent	  
 -		 val: heartbeatvalue 
 -		 event: message_sent 
 -		  
 -		  
 -----------------------------------------------------------------------------
*/

//`timescale 1 ns / 100 ps

module bench;

parameter			NUM_HOST  = 2;

// decleare dut in/out ports
	reg				clk;
	reg				rst;
	reg				connect_i;			// from app
	reg[1:0]			connect_to_host_i;		// from app

	reg				connected_i_i;			// from toe
	reg[1:0]			connected_host_addr_i_i;		// from toe
	reg[1:0]			id_i_i;				// from toe
	reg[7:0]			message_i_i;			// from toe
	reg				fifo_full_i_i;
	reg				new_message_i_i;			// will be implemented by fifo contr.

	reg				fifo_write_i_o;
	reg[7:0]			message_i_o;			// goes to fifo
	reg				end_i_o;


	reg				clk;
	reg				rst;

	reg				connected_a_i;			// from toe
	reg[1:0]			connected_host_addr_a_i;		// from toe
	reg[1:0]			id_a_i;				// from toe
	reg[7:0]			message_a_i;			// from toe
	reg				fifo_full_a_i;
	reg				new_message_a_i;			// will be implemented by fifo contr.


	reg				fifo_write_a_o;
	reg[7:0]			message_a_o;			// goes to fifo
	reg				end_a_o;


// instantiate dut
end_to_end_system dut (	  
	 	.clk,
	 	.rst,
		.id_i_i,
		.id_a_i,
	 	.connect_i,			// from app
	 	.connect_to_host_i,		// from app
	 	.connected_i_i,			// from toe
	 	.connected_host_addr_i_i,		// from toe
	 	.message_i_i,			// from toe
		.fifo_full_i_i,
		.new_message_i_i,			// will be implemented by fifo contr.

		.fifo_write_i_o,
		.message_i_o,
		.end_i_o,

	 	.clk,
	 	.rst,

	 	.connected_a_i,			// from toe
	 	.connected_host_addr_a_i,		// from toe
	 	.message_a_i,			// from toe
		.fifo_full_a_i,
		.new_message_a_i,			// will be implemented by fifo contr.

		.fifo_write_a_o,
		.message_a_o,
		.end_a_o
	);

// internal variables and events
reg	 t_fifo_write_o;
reg	 chk_connect;
reg	 t_end_o;
reg	 t1_end_o;
reg	 t2_end_o;
reg	 t3_end_o;

integer chksm_tag_done;
integer	not_done;
integer	temp;
integer statusI,statusO, mon;
reg	  start_checking;
reg	  start_checking_a;
reg [7:0] exp;
reg [7:0] exp_g;		// garbage
integer 	in,out,cfg;
integer dut_error;
integer		temp_count;
integer		temp_count_a;
integer		count_bytes;
reg		start;



//reg[499:0]	buffer_i[7:0]; 
reg[7:0]	buffer_i[499:0]; 
integer		addr_i;		// initialize to zero
integer		t1_i;
integer		temp_addr_i;

reg[7:0]	buffer_a[499:0]; 
integer		addr_a;		// initialize to zero
integer		t1_a;
integer		temp_addr_a;
reg		transfer_i2a;
reg		transfer_a2i;

event message_sent;
event reset_enable;
event reset_done;
event exit_sim;
event configure_enable;
event configure_done;
event start_initiator;
event start_acceptor;
event error;
event initiation_trigger_sent;
event waiting_for_ack_i;
event waiting_for_ack_a;
event connected_i;
event connected_a;
event comparison_done;
event handle_checksum;
event handle_time;
event handle_bodylength;
event input_stimuli_sent;
event send_message;
event transfer_message_i2a;
event transfer_message_a2i;


// clock generator
always # 1 clk = ~clk;

// dumping waveforms
initial 
begin
  	$dumpfile ("dut.vcd");
  	$dumpvars;
end

//enable if compiling with VCS
//initial 

initial begin

$vcdpluson;		 

end

// initialization
initial begin
	$display ("\n");
	$display ("################################################### \n");
//	$fdisplay (mon, "################################################### \n");
//  	$display ("STARTING SIMULATION\n");
//	$fdisplay (mon, "STARTING SIMULATION\n");
	temp			=	0;
	clk			=	'0;
    	rst			=	'0;
    	connect_i		=	'0;
	connect_to_host_i	=	'0;
    	connected_i_i		=	'0;
    	connected_a_i		=	'0;
  	connected_host_addr_i_i	=	'0;
  	connected_host_addr_a_i	=	'0;
	id_i_i			=	'0;
	id_a_i			=	'0;
	fifo_full_a_i		=	'0;
   	new_message_i_i		=	'0;
   	new_message_a_i		=	'0;
  	message_i_i		=	'0;
  	message_a_i		=	'0;
	temp_count		=	0;
	temp_count_a		=	0;
	count_bytes		=	0;
	chksm_tag_done		=	10;
	addr_i			=	0;
	addr_a			=	0;
	t1_a			=	0;
	t1_i			=	0;
	temp_addr_a		=	0;
	temp_addr_i		=	0;

  	in  = $fopen("init_out.txt","r");
  	mon = $fopen("monitor.txt","w");
	
//	$fdisplay (mon, "Initiator Name: CLIENT1 \nAcceptor Name: ORDERMATCH \n");
end

initial begin
  	#10 -> reset_enable;
  	@ (reset_done);
  	#10 -> start_initiator;
  	#1 -> start_acceptor;
end

<<<<<<< HEAD
// applying reset logic
initial
forever begin
 	@ (reset_enable);
 	@ (posedge clk)
 	$display ("Applying reset @ %0dns", $time);
   	rst = 1;
 	@ (posedge clk)
   	rst = 0;
 	$display ("Came out of Reset @ %0dns", $time);
 	-> reset_done;
end

=======
>>>>>>> f83c563eb82b7b51e483b1d7ea09393642d0a2ce
// initiate initiator  
initial 
forever begin 
	@ (start_initiator);
	@ (posedge clk)
<<<<<<< HEAD
	$display ("Initiator: Initiating a new connection @ %0dns", $time);
=======
	$display ("Initiating a new connection request @ %0dns", $time);
//	$fdisplay (mon, "Initiating a new connection requst @ %0dns", $time);
>>>>>>> f83c563eb82b7b51e483b1d7ea09393642d0a2ce
	connect_i = '1;
	connect_to_host_i  =  2'b01; 
	@ (posedge clk)
	connect_i = '0;
<<<<<<< HEAD
	-> waiting_for_ack_i;
	@connected_i;
	#7 connected_i_i = '0;
	$display ("ACK received @ %0dns", $time);

	#10000 $finish;

//	@error;
//	->exit_sim;
end

// initiate acceptor  
initial 
forever begin 
	@ (start_acceptor);
	@ (posedge clk)
	$display ("Acceptor: waiting for a new connection @ %0dns", $time);
	-> waiting_for_ack_a;
	@connected_a;
	#7 connected_a_i = '0;
	$display ("ACK received @ %0dns", $time);

//	#1000 $finish;	

//	@error;
//	->exit_sim;
end

// connection status: initiator side  
initial begin
	@(waiting_for_ack_i);
	#3 @(posedge clk)
	connected_i_i = '1;
	connected_host_addr_i_i = 2'b01;
	->connected_i;
end

// connection status: acceptor side  
initial begin
	@(waiting_for_ack_a);
	#3 @(posedge clk)
	connected_a_i = '1;
	connected_host_addr_a_i = 2'b00;
	->connected_a;
end

reg		start;

always @(*) begin

	if (fifo_write_i_o == 1 && connect_i == 0) begin
		start	=	'1;
	end else	
		start	=	'0;
end

reg[7:0]		message_temp;

always @ (posedge clk) begin

	if (start == 1) begin
		if (temp_count <1) begin
			temp_count	=	temp_count + 1;
			start_checking  = '0;
		end else begin
			buffer_i[addr_i]    = message_i_o;
			addr_i = addr_i + 1;	
			start_checking  = '1; 
		end
	end else
			start_checking	=	'0;
end


// buffer sent data from each end
always @ (posedge clk) begin

		new_message_a_i = '0;

	if (end_i_o  == 1) begin
		temp_count  = 0;
		temp_addr_i   =  addr_i;
		addr_i	 = 0;
		new_message_a_i = '1;
	end
end

always @ (*) begin
	if (t1_i == temp_addr_i-1) begin
		transfer_i2a <= '0;
		t1_i	= '0;
	end
end

always @ (posedge clk) begin

	if (new_message_a_i == 1)
		transfer_i2a <= '1;	
end

always @ (posedge clk) begin

	if (transfer_i2a == 1) begin
		message_a_i	=	buffer_i[1+t1_i];
		t1_i = t1_i + 1;
	end
end


// ------------------ acceptor -------------


reg		start_a;

always @(*) begin

	if (fifo_write_a_o == 1 ) begin
		start_a	=	'1;
	end else	
		start_a	=	'0;
end

always @ (posedge clk) begin

	if (start_a == 1) begin
		if (temp_count_a <1) begin
			temp_count_a	=	temp_count_a + 1;
			start_checking_a  = '0;
		end else begin
			buffer_a[addr_a]    = message_a_o;
			addr_a = addr_a + 1;	
			start_checking_a  = '1; 
		end
	end else
			start_checking_a	=	'0;
end


// buffer sent data from each end
always @ (posedge clk) begin

		new_message_i_i = '0;

	if (end_a_o  == 1) begin
		temp_count_a  = 0;
		temp_addr_a   =  addr_a;
		addr_a	 = 0;
		new_message_i_i = '1;
	end
end

always @ (*) begin
	if (t1_a == temp_addr_a-1) begin
		transfer_a2i <= '0;
		t1_a	= '0;
	end
end

always @ (posedge clk) begin

	if (new_message_i_i == 1)
		transfer_a2i <= '1;	
end

always @ (posedge clk) begin

	if (transfer_a2i == 1) begin
		message_i_i	=	buffer_a[1+t1_a];
		t1_a = t1_a + 1;
	end
=======
	-> waiting_for_ack;
	@connected;
	#7 connected_i = '0;
	-> input_stimuli_sent;
	$display ("ACK received from TOE: connected!! @ %0dns", $time);
//	$fdisplay (mon, "ACK received from TOE: connected!! @ %0dns", $time);
	@error;
	->exit_sim;
end

// applying reset logic
initial
forever begin
 	@ (reset_enable);
 	@ (negedge clk)
 	$display ("Applying reset @ %0dns", $time);
 //	$fdisplay (mon, "Applying reset @ %0dns", $time);
   	rst = 1;
 	@ (negedge clk)
   	rst = 0;
 //	$fdisplay (mon, "Came out of Reset @ %0dns", $time);
 	-> reset_done;
end

// send connection status
initial begin
	@(waiting_for_ack);
	#3 @(negedge clk)
	connected_i = '1;
	connected_host_addr_i = 2'b01;
	->connected;
>>>>>>> f83c563eb82b7b51e483b1d7ea09393642d0a2ce
end

endmodule


/*
// exiting simulation
initial
	@ (exit_sim)  begin

	if (dut_error == 1) begin
		$display ("Terminating simulation @ %0dns ", $time);
		$display ("SIMLUATION FAILED @ %0dns ", $time);
			$display("       Got  %h",message_o);
			$display("       Exp  %h",exp);
		$display ("################################################### \n");
	end else begin
		$display ("Terminating simulation @ %0dns ", $time);
		$display ("SIMLUATION PASSED @ %0dns ", $time);
		$display ("################################################### \n");
	end
 	#10 $finish;
end




// golden model
always @(*) begin

	chk_connect	=	connect_i;

	if (connect_i == 1) begin
		exp		= {3'b000, 1'b0, connect_to_host_i, 3'b000};	
	end


	if (fifo_write_o == 1 && connect_i == 0 ) begin
		start =  '1;
	end else 
		start = '0;
	
	t_fifo_write_o	=	fifo_write_o;
end

always @ (negedge clk) begin
	t_end_o  <= #5 end_o;

	if (t_end_o == '1)
		chksm_tag_done = 1;
end

always @ (negedge clk) begin
#4	t1_end_o  <= t_end_o;
end

always @ (posedge clk) begin

if (start == 1 ) begin
		if (temp_count <2  ) begin
			temp_count	=	temp_count + 1;
			start_checking = '0;
		end else begin
			start_checking = '1;
			if (count_bytes >= 12 && count_bytes < 15 && message_o != 8'h01) begin
				count_bytes = count_bytes + 1;
				statusO = $fscanf(in, "%h ",exp_g[7:0]);
				exp	= 8'h3b;
			end else if (count_bytes >= 39 && count_bytes < 61 && end_o != 1 && message_o != 8'h01) begin
				count_bytes = count_bytes + 1;
				statusO = $fscanf(in, "%h ",exp_g[7:0]);
				exp	= 8'h3b;
			end else if ( chksm_tag_done > 0 && chksm_tag_done <4  ) begin
				chksm_tag_done = chksm_tag_done + 1;
				statusO = $fscanf(in, "%h ",exp_g[7:0]);
				exp	= 8'h3b; 
			end else if (chksm_tag_done == 4) begin
				statusO = $fscanf(in, "%h %h ",exp[7:0], exp_g[7:0]);
				temp_count	=	0;				
				count_bytes	=	0;
				chksm_tag_done	=	0;
				-> message_sent;	
			end else begin
				count_bytes 	= 	count_bytes + 1;		// initialize at 5 
				statusO = $fscanf(in, "%h ",exp[7:0]);
			end
		end
end else
		start_checking	=	'0;
end

// jump here for comparison_done
initial
forever begin
	@ message_sent;

<<<<<<< HEAD
	repeat (2) @ (negedge clk) begin
		statusO = $fscanf(in, "%h ",exp_g[7:0]);
	end	
	
	@ (negedge clk)
=======
	#10 @ (negedge clk) 

>>>>>>> f83c563eb82b7b51e483b1d7ea09393642d0a2ce
	new_message_i = '1;
	id_i	=	2'b01;
	while (!$feof(in)) begin
      		@ (negedge clk);
		new_message_i = '0;
      		statusI = $fscanf(in,"%h ", message_i[7:0]);
		if (message_i == 8'h3b) begin
<<<<<<< HEAD
			repeat (400) @ (negedge clk);
		end
			new_message_i = '1;
	end
=======
			# 500 //-> input_stimuli_sent;
    		  		@ (negedge clk);
				new_message_i = '1;
		end
	end
			dut_error	=	'0;
			-> exit_sim;
>>>>>>> f83c563eb82b7b51e483b1d7ea09393642d0a2ce
end

always @ (posedge clk) begin
	if (start_checking) begin
		if (message_o == exp || exp == 8'h3b) begin
			$display("%0dns passed : input and output  matched",$time);
		end else begin
			dut_error	=	1;
			-> error;
		end
	end
end

endmodule

*/


/*
initial 
forever begin

	@ transfer_message_i2a;
//	@ (posedge clk);
//	while (t1_i <= temp_addr_i ) begin	
		@ (posedge clk);
		message_a_i = buffer_i[t1_i];
		t1_i = t1_i + 1;
//	end

end
*/
