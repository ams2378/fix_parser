library verilog;
use verilog.vl_types.all;
entity const is
    generic(
        supportedVersion: vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        seqResetMsg     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        logonMsg        : vl_logic_vector(0 to 7) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        logoutMsg       : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        heartBeatMsg    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        resendReqMsg    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        msgSeqH         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        garbled         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        msgSeqL         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        valid           : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        invalid         : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        unsupportedVersion: vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        invalidMsgType  : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        requiredTagMissing: vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        logon           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        heartbeat       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        resendReq       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        logout          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        reset           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        gapFill         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        business        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        possDupFlag     : integer := 13363;
        msgSeqNum       : integer := 13108;
        targetCompId    : integer := 13622;
        sourceCompId    : integer := 13369;
        beginSeqNum     : integer := 55;
        endSeqNum       : integer := 12598;
        gapFillFlag     : integer := 3224115;
        newSeqNum       : integer := 13110;
        heartbeatInt    : integer := 48;
        sendtime        : integer := 13618;
        t_beginString   : integer := 56;
        t_bodylength    : integer := 57;
        t_msgType       : integer := 13109
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of supportedVersion : constant is 1;
    attribute mti_svvh_generic_type of seqResetMsg : constant is 1;
    attribute mti_svvh_generic_type of logonMsg : constant is 1;
    attribute mti_svvh_generic_type of logoutMsg : constant is 1;
    attribute mti_svvh_generic_type of heartBeatMsg : constant is 1;
    attribute mti_svvh_generic_type of resendReqMsg : constant is 1;
    attribute mti_svvh_generic_type of msgSeqH : constant is 1;
    attribute mti_svvh_generic_type of garbled : constant is 1;
    attribute mti_svvh_generic_type of msgSeqL : constant is 1;
    attribute mti_svvh_generic_type of valid : constant is 1;
    attribute mti_svvh_generic_type of invalid : constant is 1;
    attribute mti_svvh_generic_type of unsupportedVersion : constant is 1;
    attribute mti_svvh_generic_type of invalidMsgType : constant is 1;
    attribute mti_svvh_generic_type of requiredTagMissing : constant is 1;
    attribute mti_svvh_generic_type of logon : constant is 1;
    attribute mti_svvh_generic_type of heartbeat : constant is 1;
    attribute mti_svvh_generic_type of resendReq : constant is 1;
    attribute mti_svvh_generic_type of logout : constant is 1;
    attribute mti_svvh_generic_type of reset : constant is 1;
    attribute mti_svvh_generic_type of gapFill : constant is 1;
    attribute mti_svvh_generic_type of business : constant is 1;
    attribute mti_svvh_generic_type of possDupFlag : constant is 1;
    attribute mti_svvh_generic_type of msgSeqNum : constant is 1;
    attribute mti_svvh_generic_type of targetCompId : constant is 1;
    attribute mti_svvh_generic_type of sourceCompId : constant is 1;
    attribute mti_svvh_generic_type of beginSeqNum : constant is 1;
    attribute mti_svvh_generic_type of endSeqNum : constant is 1;
    attribute mti_svvh_generic_type of gapFillFlag : constant is 1;
    attribute mti_svvh_generic_type of newSeqNum : constant is 1;
    attribute mti_svvh_generic_type of heartbeatInt : constant is 1;
    attribute mti_svvh_generic_type of sendtime : constant is 1;
    attribute mti_svvh_generic_type of t_beginString : constant is 1;
    attribute mti_svvh_generic_type of t_bodylength : constant is 1;
    attribute mti_svvh_generic_type of t_msgType : constant is 1;
end const;
