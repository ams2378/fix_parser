module tagsort (




);





