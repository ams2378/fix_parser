library verilog;
use verilog.vl_types.all;
entity parser_test is
end parser_test;
