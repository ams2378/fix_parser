library verilog;
use verilog.vl_types.all;
entity fix_engine_test is
end fix_engine_test;
