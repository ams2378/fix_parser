
`ifndef _my_incl_vh_
`define _my_incl_vh_

`define logon 1 //3'b001;
`define business 7 // 3'b111;
`define logout 4 //3'b100;
`define heartbeat 2 //3'b010;


`endif
